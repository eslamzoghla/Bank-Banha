module Rom(addr,wtime);
  // -------------------------- Inputs Declarations ---------------------------- //
  input [4:0]addr;
  // -------------------------- Outputs Declarations ---------------------------- // 
  output [4:0]wtime;
  // -------------------------- Reg Declarations ---------------------------- //
  reg [4:0]  rom [0:31];
  // ----------------------- Sequential  Logic  -------------------------------- //
  always@(*)
  begin //<<<<<<<<<<<<<<<<<<<<<<<<<<<< Start Always block >>>>>>>>>>>>>>>>>>>>>>>>>>
    case(addr)
	 
    //(1 teller)  
    5'b01000 : rom[addr]<=5'b00000;//0
    5'b01001 : rom[addr]<=5'b00011;//3
    5'b01010 : rom[addr]<=5'b00110;//6
    5'b01011 : rom[addr]<=5'b01001;//9
    5'b01100 : rom[addr]<=5'b01100;//12
    5'b01101 : rom[addr]<=5'b01111;//15
    5'b01110 : rom[addr]<=5'b10010;//18
    5'b01111 : rom[addr]<=5'b10101;//21
    
    //(2 tellers)
    5'b10000 : rom[addr]<=5'b00000;//0
    5'b10001 : rom[addr]<=5'b00011;//3
    5'b10010 : rom[addr]<=5'b00101;//5
    5'b10011 : rom[addr]<=5'b00110;//6
    5'b10100 : rom[addr]<=5'b01000;//8
    5'b10101 : rom[addr]<=5'b01001;//9
    5'b10110 : rom[addr]<=5'b01011;//11
    5'b10111 : rom[addr]<=5'b01100;//12
    
    //(3 tellers)
    5'b11000 : rom[addr]<=5'b00000;//0
    5'b11001 : rom[addr]<=5'b00011;//3
    5'b11010 : rom[addr]<=5'b00100;//4
    5'b11011 : rom[addr]<=5'b00101;//5
    5'b11100 : rom[addr]<=5'b00110;//6
    5'b11101 : rom[addr]<=5'b00111;//7
    5'b11110 : rom[addr]<=5'b01000;//8
    5'b11111 : rom[addr]<=5'b01001;//9
    
    default : rom[addr]<=5'b00000;//0
   endcase  
  end//<<<<<<<<<<<<<<<<<<<<<<<<<<<< End Always block >>>>>>>>>>>>>>>>>>>>>>>>>>
  
      assign wtime =rom[addr];
  
endmodule

	// ----------------------------- End of File --------------------------------- //
	// --------------------------------------------------------------------------- //
